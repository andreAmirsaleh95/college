module memReg(); 
endmodule
